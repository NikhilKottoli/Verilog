`timescale 1ns/1ns
`include "Hello.v"

module testbase;
    reg W,X,Y,Z;
    wire A,B,C,D;
    gate output
endmodule